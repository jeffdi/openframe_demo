magic
tech sky130A
magscale 1 2
timestamp 1686347941
<< nwell >>
rect 1066 56837 58918 57403
rect 1066 55749 58918 56315
rect 1066 54661 58918 55227
rect 1066 53573 58918 54139
rect 1066 52485 58918 53051
rect 1066 51397 58918 51963
rect 1066 50309 58918 50875
rect 1066 49221 58918 49787
rect 1066 48133 58918 48699
rect 1066 47045 58918 47611
rect 1066 45957 58918 46523
rect 1066 44869 58918 45435
rect 1066 43781 58918 44347
rect 1066 42693 58918 43259
rect 1066 41605 58918 42171
rect 1066 40517 58918 41083
rect 1066 39429 58918 39995
rect 1066 38341 58918 38907
rect 1066 37253 58918 37819
rect 1066 36165 58918 36731
rect 1066 35077 58918 35643
rect 1066 33989 58918 34555
rect 1066 32901 58918 33467
rect 1066 31813 58918 32379
rect 1066 30725 58918 31291
rect 1066 29637 58918 30203
rect 1066 28549 58918 29115
rect 1066 27461 58918 28027
rect 1066 26373 58918 26939
rect 1066 25285 58918 25851
rect 1066 24197 58918 24763
rect 1066 23109 58918 23675
rect 1066 22021 58918 22587
rect 1066 20933 58918 21499
rect 1066 19845 58918 20411
rect 1066 18757 58918 19323
rect 1066 17669 58918 18235
rect 1066 16581 58918 17147
rect 1066 15493 58918 16059
rect 1066 14405 58918 14971
rect 1066 13317 58918 13883
rect 1066 12229 58918 12795
rect 1066 11141 58918 11707
rect 1066 10053 58918 10619
rect 1066 8965 58918 9531
rect 1066 7877 58918 8443
rect 1066 6789 58918 7355
rect 1066 5701 58918 6267
rect 1066 4613 58918 5179
rect 1066 3525 58918 4091
rect 1066 2437 58918 3003
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 1104 2128 58880 57712
<< metal2 >>
rect 3974 59200 4030 60000
rect 4434 59200 4490 60000
rect 4894 59200 4950 60000
rect 5354 59200 5410 60000
rect 5814 59200 5870 60000
rect 6274 59200 6330 60000
rect 6734 59200 6790 60000
rect 7194 59200 7250 60000
rect 7654 59200 7710 60000
rect 8114 59200 8170 60000
rect 8574 59200 8630 60000
rect 9034 59200 9090 60000
rect 9494 59200 9550 60000
rect 9954 59200 10010 60000
rect 10414 59200 10470 60000
rect 10874 59200 10930 60000
rect 11334 59200 11390 60000
rect 11794 59200 11850 60000
rect 12254 59200 12310 60000
rect 12714 59200 12770 60000
rect 13174 59200 13230 60000
rect 13634 59200 13690 60000
rect 14094 59200 14150 60000
rect 14554 59200 14610 60000
rect 15014 59200 15070 60000
rect 15474 59200 15530 60000
rect 15934 59200 15990 60000
rect 16394 59200 16450 60000
rect 16854 59200 16910 60000
rect 17314 59200 17370 60000
rect 17774 59200 17830 60000
rect 18234 59200 18290 60000
rect 18694 59200 18750 60000
rect 19154 59200 19210 60000
rect 19614 59200 19670 60000
rect 20074 59200 20130 60000
rect 20534 59200 20590 60000
rect 20994 59200 21050 60000
rect 21454 59200 21510 60000
rect 21914 59200 21970 60000
rect 22374 59200 22430 60000
rect 22834 59200 22890 60000
rect 23294 59200 23350 60000
rect 23754 59200 23810 60000
rect 24214 59200 24270 60000
rect 24674 59200 24730 60000
rect 25134 59200 25190 60000
rect 25594 59200 25650 60000
rect 26054 59200 26110 60000
rect 26514 59200 26570 60000
rect 26974 59200 27030 60000
rect 27434 59200 27490 60000
rect 27894 59200 27950 60000
rect 28354 59200 28410 60000
rect 28814 59200 28870 60000
rect 29274 59200 29330 60000
rect 29734 59200 29790 60000
rect 30194 59200 30250 60000
rect 30654 59200 30710 60000
rect 31114 59200 31170 60000
rect 31574 59200 31630 60000
rect 32034 59200 32090 60000
rect 32494 59200 32550 60000
rect 32954 59200 33010 60000
rect 33414 59200 33470 60000
rect 33874 59200 33930 60000
rect 34334 59200 34390 60000
rect 34794 59200 34850 60000
rect 35254 59200 35310 60000
rect 35714 59200 35770 60000
rect 36174 59200 36230 60000
rect 36634 59200 36690 60000
rect 37094 59200 37150 60000
rect 37554 59200 37610 60000
rect 38014 59200 38070 60000
rect 38474 59200 38530 60000
rect 38934 59200 38990 60000
rect 39394 59200 39450 60000
rect 39854 59200 39910 60000
rect 40314 59200 40370 60000
rect 40774 59200 40830 60000
rect 41234 59200 41290 60000
rect 41694 59200 41750 60000
rect 42154 59200 42210 60000
rect 42614 59200 42670 60000
rect 43074 59200 43130 60000
rect 43534 59200 43590 60000
rect 43994 59200 44050 60000
rect 44454 59200 44510 60000
rect 44914 59200 44970 60000
rect 45374 59200 45430 60000
rect 45834 59200 45890 60000
rect 46294 59200 46350 60000
rect 46754 59200 46810 60000
rect 47214 59200 47270 60000
rect 47674 59200 47730 60000
rect 48134 59200 48190 60000
rect 48594 59200 48650 60000
rect 49054 59200 49110 60000
rect 49514 59200 49570 60000
rect 49974 59200 50030 60000
rect 50434 59200 50490 60000
rect 50894 59200 50950 60000
rect 51354 59200 51410 60000
rect 51814 59200 51870 60000
rect 52274 59200 52330 60000
rect 52734 59200 52790 60000
rect 53194 59200 53250 60000
rect 53654 59200 53710 60000
rect 54114 59200 54170 60000
rect 54574 59200 54630 60000
rect 55034 59200 55090 60000
rect 55494 59200 55550 60000
rect 55954 59200 56010 60000
<< obsm2 >>
rect 4214 59144 4378 59200
rect 4546 59144 4838 59200
rect 5006 59144 5298 59200
rect 5466 59144 5758 59200
rect 5926 59144 6218 59200
rect 6386 59144 6678 59200
rect 6846 59144 7138 59200
rect 7306 59144 7598 59200
rect 7766 59144 8058 59200
rect 8226 59144 8518 59200
rect 8686 59144 8978 59200
rect 9146 59144 9438 59200
rect 9606 59144 9898 59200
rect 10066 59144 10358 59200
rect 10526 59144 10818 59200
rect 10986 59144 11278 59200
rect 11446 59144 11738 59200
rect 11906 59144 12198 59200
rect 12366 59144 12658 59200
rect 12826 59144 13118 59200
rect 13286 59144 13578 59200
rect 13746 59144 14038 59200
rect 14206 59144 14498 59200
rect 14666 59144 14958 59200
rect 15126 59144 15418 59200
rect 15586 59144 15878 59200
rect 16046 59144 16338 59200
rect 16506 59144 16798 59200
rect 16966 59144 17258 59200
rect 17426 59144 17718 59200
rect 17886 59144 18178 59200
rect 18346 59144 18638 59200
rect 18806 59144 19098 59200
rect 19266 59144 19558 59200
rect 19726 59144 20018 59200
rect 20186 59144 20478 59200
rect 20646 59144 20938 59200
rect 21106 59144 21398 59200
rect 21566 59144 21858 59200
rect 22026 59144 22318 59200
rect 22486 59144 22778 59200
rect 22946 59144 23238 59200
rect 23406 59144 23698 59200
rect 23866 59144 24158 59200
rect 24326 59144 24618 59200
rect 24786 59144 25078 59200
rect 25246 59144 25538 59200
rect 25706 59144 25998 59200
rect 26166 59144 26458 59200
rect 26626 59144 26918 59200
rect 27086 59144 27378 59200
rect 27546 59144 27838 59200
rect 28006 59144 28298 59200
rect 28466 59144 28758 59200
rect 28926 59144 29218 59200
rect 29386 59144 29678 59200
rect 29846 59144 30138 59200
rect 30306 59144 30598 59200
rect 30766 59144 31058 59200
rect 31226 59144 31518 59200
rect 31686 59144 31978 59200
rect 32146 59144 32438 59200
rect 32606 59144 32898 59200
rect 33066 59144 33358 59200
rect 33526 59144 33818 59200
rect 33986 59144 34278 59200
rect 34446 59144 34738 59200
rect 34906 59144 35198 59200
rect 35366 59144 35658 59200
rect 35826 59144 36118 59200
rect 36286 59144 36578 59200
rect 36746 59144 37038 59200
rect 37206 59144 37498 59200
rect 37666 59144 37958 59200
rect 38126 59144 38418 59200
rect 38586 59144 38878 59200
rect 39046 59144 39338 59200
rect 39506 59144 39798 59200
rect 39966 59144 40258 59200
rect 40426 59144 40718 59200
rect 40886 59144 41178 59200
rect 41346 59144 41638 59200
rect 41806 59144 42098 59200
rect 42266 59144 42558 59200
rect 42726 59144 43018 59200
rect 43186 59144 43478 59200
rect 43646 59144 43938 59200
rect 44106 59144 44398 59200
rect 44566 59144 44858 59200
rect 45026 59144 45318 59200
rect 45486 59144 45778 59200
rect 45946 59144 46238 59200
rect 46406 59144 46698 59200
rect 46866 59144 47158 59200
rect 47326 59144 47618 59200
rect 47786 59144 48078 59200
rect 48246 59144 48538 59200
rect 48706 59144 48998 59200
rect 49166 59144 49458 59200
rect 49626 59144 49918 59200
rect 50086 59144 50378 59200
rect 50546 59144 50838 59200
rect 51006 59144 51298 59200
rect 51466 59144 51758 59200
rect 51926 59144 52218 59200
rect 52386 59144 52678 59200
rect 52846 59144 53138 59200
rect 53306 59144 53598 59200
rect 53766 59144 54058 59200
rect 54226 59144 54518 59200
rect 54686 59144 54978 59200
rect 55146 59144 55438 59200
rect 55606 59144 55898 59200
rect 4214 2139 56008 59144
<< obsm3 >>
rect 4210 2143 50606 57697
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< labels >>
rlabel metal2 s 3974 59200 4030 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 17774 59200 17830 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 19154 59200 19210 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 20534 59200 20590 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 21914 59200 21970 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 23294 59200 23350 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 24674 59200 24730 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 26054 59200 26110 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 27434 59200 27490 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 28814 59200 28870 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 30194 59200 30250 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5354 59200 5410 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 31574 59200 31630 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 32954 59200 33010 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 34334 59200 34390 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 35714 59200 35770 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 37094 59200 37150 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 38474 59200 38530 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 39854 59200 39910 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 41234 59200 41290 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 42614 59200 42670 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 43994 59200 44050 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 6734 59200 6790 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 45374 59200 45430 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 46754 59200 46810 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 48134 59200 48190 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 49514 59200 49570 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 50894 59200 50950 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 52274 59200 52330 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 53654 59200 53710 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 55034 59200 55090 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8114 59200 8170 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 9494 59200 9550 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 10874 59200 10930 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 12254 59200 12310 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 13634 59200 13690 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 15014 59200 15070 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 16394 59200 16450 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4434 59200 4490 60000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 18234 59200 18290 60000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 19614 59200 19670 60000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 20994 59200 21050 60000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 22374 59200 22430 60000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 23754 59200 23810 60000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 25134 59200 25190 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 26514 59200 26570 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 27894 59200 27950 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 29274 59200 29330 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 30654 59200 30710 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 5814 59200 5870 60000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 32034 59200 32090 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 33414 59200 33470 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 34794 59200 34850 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 36174 59200 36230 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 37554 59200 37610 60000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 38934 59200 38990 60000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 40314 59200 40370 60000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 41694 59200 41750 60000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 43074 59200 43130 60000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 44454 59200 44510 60000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 7194 59200 7250 60000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 45834 59200 45890 60000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 47214 59200 47270 60000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 48594 59200 48650 60000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 49974 59200 50030 60000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 51354 59200 51410 60000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 52734 59200 52790 60000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 54114 59200 54170 60000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 55494 59200 55550 60000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 8574 59200 8630 60000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 9954 59200 10010 60000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 11334 59200 11390 60000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 12714 59200 12770 60000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 14094 59200 14150 60000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 15474 59200 15530 60000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 16854 59200 16910 60000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4894 59200 4950 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 18694 59200 18750 60000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 20074 59200 20130 60000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 21454 59200 21510 60000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 22834 59200 22890 60000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 24214 59200 24270 60000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 25594 59200 25650 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 26974 59200 27030 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 28354 59200 28410 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 29734 59200 29790 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 31114 59200 31170 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 6274 59200 6330 60000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 32494 59200 32550 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 33874 59200 33930 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 35254 59200 35310 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 36634 59200 36690 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 38014 59200 38070 60000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 39394 59200 39450 60000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 40774 59200 40830 60000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 42154 59200 42210 60000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 43534 59200 43590 60000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 44914 59200 44970 60000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7654 59200 7710 60000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 46294 59200 46350 60000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 47674 59200 47730 60000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 49054 59200 49110 60000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 50434 59200 50490 60000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 51814 59200 51870 60000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 53194 59200 53250 60000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 54574 59200 54630 60000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 55954 59200 56010 60000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9034 59200 9090 60000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 10414 59200 10470 60000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 11794 59200 11850 60000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 13174 59200 13230 60000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 14554 59200 14610 60000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 15934 59200 15990 60000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 17314 59200 17370 60000 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1200844
string GDS_FILE /home/jeffdi/openframe_demo/openlane/user_proj_example/runs/23_06_09_14_57/results/signoff/user_proj_example.magic.gds
string GDS_START 167052
<< end >>

